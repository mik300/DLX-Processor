LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;
--USE IEEE.numeric_std.all;
--USE WORK.CONSTANTS.ALL;

ENTITY DRAM IS
	GENERIC( ADDR_LEN : NATURAL;
			 DATA_LEN : NATURAL);
	PORT (CLK:      IN  std_logic;
          RESET: 	IN  std_logic;
	      WR: 		IN  std_logic;
	      ADDRESS:	IN  std_logic_vector(ADDR_LEN-1 DOWNTO 0);
	      DATAIN: 	IN  std_logic_vector(DATA_LEN-1 DOWNTO 0); --1 WRITE AT A TIME
          DATAOUT:  OUT std_logic_vector(DATA_LEN-1 DOWNTO 0));

END DRAM;

ARCHITECTURE A OF DRAM IS

    -- suggested structures
	SUBTYPE REG_ADDR IS NATURAL RANGE 0 TO 2**ADDR_LEN -1; -- using natural type -- 2**ADDR_LEN Registers
	TYPE REG_ARRAY IS ARRAY(REG_ADDR) OF STD_LOGIC_VECTOR(DATA_LEN-1 DOWNTO 0);  --Each row has DATA_LEN bits
	SIGNAL REGISTERS: REG_ARRAY := (OTHERS => (OTHERS => '0'));

BEGIN

	--REGISTERS(0) <= x"00000000";

	WRITE :  PROCESS(CLK, RESET) 
	BEGIN 
		IF (RESET = '1') THEN
			REGISTERS <= (OTHERS => (OTHERS => '0'));
		ELSIF (RISING_EDGE(CLK)) THEN
			IF(WR = '1') THEN 
				REGISTERS(CONV_INTEGER(ADDRESS)) <= DATAIN; 
			END IF;
		END IF;
	END PROCESS WRITE;

	Read1 : PROCESS(ADDRESS, REGISTERS) 
	BEGIN
		DATAOUT <= REGISTERS(CONV_INTEGER(ADDRESS));				
	END PROCESS Read1;


END A;

CONFIGURATION CFG_RF_BEH OF DRAM IS
  FOR A
  END FOR;
END CONFIGURATION;
