!<symlink>��/ e d a / d k / n a n g a t e 4 5 / l e f / N a n g a t e O p e n C e l l L i b r a r y . l e f   